// Plik zawieraj�cy definicje do timingu vga wed�ug standardu VESA

`ifndef _vesa_vga_vh_
`define _vesa_vga_vh

`define VS_START 601
`define VS_DURATION 4
`define VS_END 605

`define HS_START 840
`define HS_DURATION 128
`define HS_END 968

`define HB_START 800
`define HB_DURATION 255
`define HB_END 1055

`define VB_START 600
`define VB_DURATION 27
`define VB_END 627

`define VC_MAX 627
`define HC_MAX 1055

`endif